package test_pkg;

    // Конфигурация тестового сценария

    `include "cfg.sv"  

    // Пакет

    `include "packet.sv"

    // Генератор

    `include "gen.sv"

    // Драйвер

    `include "driver.sv"

    // Монитор

    `include "monitor.sv"

    // Агент

    `include "agent.sv"

endpackage