class env_base;
    
    master_data_aligner_agent_base master;
    slave_data_aligner_agent_base  slave;
    checker_data_aligner_base      check;

    function new();
        master  = new();
        slave   = new();
        check   = new();
    endfunction

    virtual task run();
        fork
            master.run();
            slave .run();
            check .run();
        join
    endtask
    
endclass