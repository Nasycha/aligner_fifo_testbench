package test_pkg;

    // Конфигурация тестового сценария

    `include "data_align_cfg.sv"  

    // Пакет

    `include "data_align_packet.sv"

    // Генератор

    `include "data_align_gen.sv"

    // Драйвер

    `include "data_align_driver.sv"

    // Монитор

    `include "data_align_monitor.sv"

    // Агент

    `include "data_align_agent.sv"

    // Проверка

    `include "data_align_checker.sv"

    // Окружение

    `include "data_align_env.sv"

    // Тест

    `include "data_align_test.sv"

endpackage